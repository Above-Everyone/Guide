module src

// test := {
//   "username": "Webhook",
//   "avatar_url": "https://i.imgur.com/4M34hi2.png",
//   "content": "Text message. Up to 2000 characters.",
//   "embeds": [
//     {
//       "author": {
//         "name": "Birdie♫",
//         "url": "https://www.reddit.com/r/cats/",
//         "icon_url": "https://i.imgur.com/R66g1Pe.jpg"
//       },
//       "title": "Title",
//       "url": "https://google.com/",
//       "description": "Text message. You can use Markdown here. *Italic* **bold** __underline__ ~~strikeout~~ [hyperlink](https://google.com) `code`",
//       "color": 15258703,
//       "fields": [
//         {
//           "name": "Application",
//           "value": "{YM_APPLICATION_TYPE}",
//           "inline": true
//         },
//         {
//           "name": "IP Address",
//           "value": "{CLIENTS_IP_ADDRESS}",
//           "inline": true
//         },
//         {
//           "name": "Item Search Query",
//           "value": "{CLIENTS_SEARCH_QUERY}",
// 		  "inline": true
//         },
//         {
//          "name": "Results Type",
//           "value": "{YM_RESULT_TYPE}",
// 		  "inline": true
//         },
//         {
//          "name": "Results Count",
//           "value": "{YM_RESULT_COUNT}",
// 		  "inline": true
//         },
//         {
//          "name": "Current Time",
//           "value": "{CURRENT_TIME}",
// 		  "inline": true
//         }
//       ],
//       "thumbnail": {
//         "url": "https://upload.wikimedia.org/wikipedia/commons/3/38/4-Nature-Wallpapers-2014-1_ukaavUI.jpg"
//       },
//       "image": {
//         "url": "https://upload.wikimedia.org/wikipedia/commons/5/5a/A_picture_from_China_every_day_108.jpg"
//       },
//       "footer": {
//         "text": "Woah! So cool! :smirk:",
//         "icon_url": "https://i.imgur.com/fKL31aD.jpg"
//       }
//     }
//   ]
// }