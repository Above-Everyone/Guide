module db

pub struct WTB 
{
	pub mut:
		posted_timestamp	string
		wtb_price			string
		item				Item
}